module hexa (
		output wire [6:0] seg1, seg2, seg3, seg4, seg5, seg6,
		output wire [7:0] leds,
		input wire [31:0] binary
);

assign seg1 = (binary[3:0] == 4'b0000) ? 7'b1000000 : // 0
              (binary[3:0] == 4'b0001) ? 7'b1111001 : // 1
              (binary[3:0] == 4'b0010) ? 7'b0100100 : // 2
              (binary[3:0] == 4'b0011) ? 7'b0110000 : // 3
              (binary[3:0] == 4'b0100) ? 7'b0011001 : // 4
              (binary[3:0] == 4'b0101) ? 7'b0010010 : // 5
              (binary[3:0] == 4'b0110) ? 7'b0000010 : // 6
              (binary[3:0] == 4'b0111) ? 7'b1111000 : // 7
              (binary[3:0] == 4'b1000) ? 7'b0000000 : // 8
              (binary[3:0] == 4'b1001) ? 7'b0010000 : // 9
              (binary[3:0] == 4'b1010) ? 7'b0001000 : // A
              (binary[3:0] == 4'b1011) ? 7'b0000011 : // b
              (binary[3:0] == 4'b1100) ? 7'b1000110 : // C
              (binary[3:0] == 4'b1101) ? 7'b0100001 : // d
              (binary[3:0] == 4'b1110) ? 7'b0000110 : // E
              (binary[3:0] == 4'b1111) ? 7'b0001110 : // F
                                         7'b1111111 ; // off

assign seg2 = (binary[7:4] == 4'b0000) ? 7'b1000000 : // 0
              (binary[7:4] == 4'b0001) ? 7'b1111001 : // 1
              (binary[7:4] == 4'b0010) ? 7'b0100100 : // 2
              (binary[7:4] == 4'b0011) ? 7'b0110000 : // 3
              (binary[7:4] == 4'b0100) ? 7'b0011001 : // 4
              (binary[7:4] == 4'b0101) ? 7'b0010010 : // 5
              (binary[7:4] == 4'b0110) ? 7'b0000010 : // 6
              (binary[7:4] == 4'b0111) ? 7'b1111000 : // 7
              (binary[7:4] == 4'b1000) ? 7'b0000000 : // 8
              (binary[7:4] == 4'b1001) ? 7'b0010000 : // 9
              (binary[7:4] == 4'b1010) ? 7'b0001000 : // A
              (binary[7:4] == 4'b1011) ? 7'b0000011 : // b
              (binary[7:4] == 4'b1100) ? 7'b1000110 : // C
              (binary[7:4] == 4'b1101) ? 7'b0100001 : // d
              (binary[7:4] == 4'b1110) ? 7'b0000110 : // E
              (binary[7:4] == 4'b1111) ? 7'b0001110 : // F
                                         7'b1111111 ; // off

assign seg3 = (binary[11:8] == 4'b0000) ? 7'b1000000 : // 0
              (binary[11:8] == 4'b0001) ? 7'b1111001 : // 1
              (binary[11:8] == 4'b0010) ? 7'b0100100 : // 2
              (binary[11:8] == 4'b0011) ? 7'b0110000 : // 3
              (binary[11:8] == 4'b0100) ? 7'b0011001 : // 4
              (binary[11:8] == 4'b0101) ? 7'b0010010 : // 5
              (binary[11:8] == 4'b0110) ? 7'b0000010 : // 6
              (binary[11:8] == 4'b0111) ? 7'b1111000 : // 7
              (binary[11:8] == 4'b1000) ? 7'b0000000 : // 8
              (binary[11:8] == 4'b1001) ? 7'b0010000 : // 9
              (binary[11:8] == 4'b1010) ? 7'b0001000 : // A
              (binary[11:8] == 4'b1011) ? 7'b0000011 : // b
              (binary[11:8] == 4'b1100) ? 7'b1000110 : // C
              (binary[11:8] == 4'b1101) ? 7'b0100001 : // d
              (binary[11:8] == 4'b1110) ? 7'b0000110 : // E
              (binary[11:8] == 4'b1111) ? 7'b0001110 : // F
                                         7'b1111111 ; // off
													  
assign seg4 = (binary[15:12] == 4'b0000) ? 7'b1000000 : // 0
              (binary[15:12] == 4'b0001) ? 7'b1111001 : // 1
              (binary[15:12] == 4'b0010) ? 7'b0100100 : // 2
              (binary[15:12] == 4'b0011) ? 7'b0110000 : // 3
              (binary[15:12] == 4'b0100) ? 7'b0011001 : // 4
              (binary[15:12] == 4'b0101) ? 7'b0010010 : // 5
              (binary[15:12] == 4'b0110) ? 7'b0000010 : // 6
              (binary[15:12] == 4'b0111) ? 7'b1111000 : // 7
              (binary[15:12] == 4'b1000) ? 7'b0000000 : // 8
              (binary[15:12] == 4'b1001) ? 7'b0010000 : // 9
              (binary[15:12] == 4'b1010) ? 7'b0001000 : // A
              (binary[15:12] == 4'b1011) ? 7'b0000011 : // b
              (binary[15:12] == 4'b1100) ? 7'b1000110 : // C
              (binary[15:12] == 4'b1101) ? 7'b0100001 : // d
              (binary[15:12] == 4'b1110) ? 7'b0000110 : // E
              (binary[15:12] == 4'b1111) ? 7'b0001110 : // F
                                         7'b1111111 ; // off
													  
assign seg5 = (binary[19:16] == 4'b0000) ? 7'b1000000 : // 0
              (binary[19:16] == 4'b0001) ? 7'b1111001 : // 1
              (binary[19:16] == 4'b0010) ? 7'b0100100 : // 2
              (binary[19:16] == 4'b0011) ? 7'b0110000 : // 3
              (binary[19:16] == 4'b0100) ? 7'b0011001 : // 4
              (binary[19:16] == 4'b0101) ? 7'b0010010 : // 5
              (binary[19:16] == 4'b0110) ? 7'b0000010 : // 6
              (binary[19:16] == 4'b0111) ? 7'b1111000 : // 7
              (binary[19:16] == 4'b1000) ? 7'b0000000 : // 8
              (binary[19:16] == 4'b1001) ? 7'b0010000 : // 9
              (binary[19:16] == 4'b1010) ? 7'b0001000 : // A
              (binary[19:16] == 4'b1011) ? 7'b0000011 : // b
              (binary[19:16] == 4'b1100) ? 7'b1000110 : // C
              (binary[19:16] == 4'b1101) ? 7'b0100001 : // d
              (binary[19:16] == 4'b1110) ? 7'b0000110 : // E
              (binary[19:16] == 4'b1111) ? 7'b0001110 : // F
                                         7'b1111111 ; // off
													  
assign seg6 = (binary[23:20] == 4'b0000) ? 7'b1000000 : // 0
              (binary[23:20] == 4'b0001) ? 7'b1111001 : // 1
              (binary[23:20] == 4'b0010) ? 7'b0100100 : // 2
              (binary[23:20] == 4'b0011) ? 7'b0110000 : // 3
              (binary[23:20] == 4'b0100) ? 7'b0011001 : // 4
              (binary[23:20] == 4'b0101) ? 7'b0010010 : // 5
              (binary[23:20] == 4'b0110) ? 7'b0000010 : // 6
              (binary[23:20] == 4'b0111) ? 7'b1111000 : // 7
              (binary[23:20] == 4'b1000) ? 7'b0000000 : // 8
              (binary[23:20] == 4'b1001) ? 7'b0010000 : // 9
              (binary[23:20] == 4'b1010) ? 7'b0001000 : // A
              (binary[23:20] == 4'b1011) ? 7'b0000011 : // b
              (binary[23:20] == 4'b1100) ? 7'b1000110 : // C
              (binary[23:20] == 4'b1101) ? 7'b0100001 : // d
              (binary[23:20] == 4'b1110) ? 7'b0000110 : // E
              (binary[23:20] == 4'b1111) ? 7'b0001110 : // F
                                         7'b1111111 ; // off
			
assign leds = binary[31:24];
													  
endmodule